library IEEE;
use IEEE.STD_LOGIC_1164.ALL;

--nothing special. just common i2c slowdown
entity slower is
	generic (                                          
	SDA_SLOW_BITS 	: STD_LOGIC_VECTOR(0 to 271) := b"10011111111111100000000000000000000111111111111110000000011111111000011111111110000000000000000000011110000000011111100001111000000001111111111110000111111000000000000000011110000000000001111111111000000000000000000000000000011111100000000000000000000000011111111111111001";
   SDA_FAST_BITS 	: STD_LOGIC_VECTOR(0 to 271) := b"10011111111111100000000000000000000111111111111110000000011111111000011111111110000000000000000000011110000000011111100001111000000001111111111110000111111111100000000000000000000000000001111110000000000000000111111110000000011111100000000000000000000000011110000111111001";
   SCL_BITS 		: STD_LOGIC_VECTOR(0 to 271) := b"11001100110011001100110011001100110011000011001100110011001100110011001100110000110011001100110011001100110011001100001100110011001100110011001100110011000011001100110011001100110011001100110000110011001100110011001100110011001100001100110011001100110011001100110011000011"
  );
    Port ( CLK3 : in  STD_LOGIC;
           to_slow : in  STD_LOGIC;
			  to_do: in STD_LOGIC;
           SCL : out  STD_LOGIC := '1';
           SDA : out  STD_LOGIC := '1');
end slower;

architecture arch of slower is
signal p_do: STD_LOGIC := '0';
signal i2ccnt: integer range 0 to 271 := 271;
begin

process(CLK3, i2ccnt) is
begin
	if rising_edge(CLK3) then
		if i2ccnt /= 271 then
			i2ccnt <= i2ccnt + 1;
		else
			if p_do /= to_do then
				p_do <= to_do;
				i2ccnt <= 0;
			end if;
		end if;
	end if;
	
	if ((to_slow = '1') and (SDA_SLOW_BITS(i2ccnt) = '1')) or ((to_slow = '0') and (SDA_FAST_BITS(i2ccnt) = '1')) then
		SDA <= 'Z';
	else
		SDA <= '0';
	end if;
		
	if SCL_BITS(i2ccnt) = '1' then
		SCL <= 'Z';
	else
		SCL <= '0';
	end if;
    
  end process;

end arch;

